module Counter();

endmodule // Counter