module StateMachine();
endmodule
